module adder #(
    parameter CLK_HZ = 25_000_000,
    parameter DEBOUNCE_MS = 10,
    parameter ACTIVE_LOW = 0,
    parameter MAX_DATA = 16,
    parameter WIDTH = $clog2(MAX_DATA)
) (
    input clk_25mhz,
    input [3:0] btn,
    output logic [WIDTH-1:0] led
);

  logic [2:0] btn_pressed;

  debounce #(
      .CLK_HZ(CLK_HZ),
      .DEBOUNCE_MS(DEBOUNCE_MS),
      .ACTIVE_LOW(ACTIVE_LOW)
  ) debounce_u0 (
      .clk(clk_25mhz),
      .btn_i(btn[0]),
      .pressed(btn_pressed[0])
  );

  debounce #(
      .CLK_HZ(CLK_HZ),
      .DEBOUNCE_MS(DEBOUNCE_MS),
      .ACTIVE_LOW(ACTIVE_LOW)
  ) debounce_u1 (
      .clk(clk_25mhz),
      .btn_i(btn[1]),
      .pressed(btn_pressed[1])
  );

  debounce #(
      .CLK_HZ(CLK_HZ),
      .DEBOUNCE_MS(DEBOUNCE_MS),
      .ACTIVE_LOW(ACTIVE_LOW)
  ) debounce_u2 (
      .clk(clk_25mhz),
      .btn_i(btn[2]),
      .pressed(btn_pressed[2])
  );

  always_ff @(posedge clk_25mhz) begin
    if (btn_pressed[0]) begin
        led <= led + 1;
    end else if (btn_pressed[1]) begin
        led <= led + (1 << 1);
    end else if (btn_pressed[2]) begin
        led <= led + (1 << 2);
    end else begin
        led <= led;
    end
  end

endmodule
